///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: pwm.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::SmartFusion> <Die::A2F200M3F> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 
`timescale <time_units> / <precision>

module pwm( clk, duty_cycle, period, pwm_out );
input port1, port2;
output port3;
inout port4;

<statements>

endmodule

