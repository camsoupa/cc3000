`timescale 1ns/1ns

module testbench();

localparam APB_DWIDTH = 32;

reg  SYSCLK;      
reg  SYSRSTN;     
wire PCLK;        
wire PRESETN;     
wire [31:0] PADDR;      
wire PENABLE;     
wire PWRITE;      
wire [APB_DWIDTH-1:0] PWDATA;     
wire [APB_DWIDTH-1:0] PRDATA;     
wire [APB_DWIDTH-1:0] PRDATA_0;     
wire [APB_DWIDTH-1:0] PRDATA_1;     
wire [15:0] PSEL;
         
wire [255:0] INTERRUPT;   
wire [31:0]  GP_OUT;      
wire [31:0]  GP_IN;       
wire FINISHED;  
wire FAILED;

wire Logic0 = 1'b0;
wire Logic1 = 1'b1;    


// ********************************************************************************
// Clocks and Reset


initial
 begin
  SYSRSTN <= 1'b0;
  #100;
  SYSRSTN <= 1'b1;
 end

// Clock is 100MHz
always
 begin
   SYSCLK <= 1'b0;
   #5;
   SYSCLK <= 1'b1;
   #5;
 end
 
   
// ********************************************************************************
// APB Master  

BFM_APB  #(.VECTFILE     ("user_tb.vec") )
     UBFM (.SYSCLK       (SYSCLK), 
           .SYSRSTN      (SYSRSTN), 
           .PCLK         (PCLK), 
           .PRESETN      (PRESETN), 
           .PADDR        (PADDR), 
           .PENABLE      (PENABLE), 
           .PWRITE       (PWRITE), 
           .PWDATA       (PWDATA), 
           .PRDATA       (PRDATA), 
           .PREADY       (Logic1), 
           .PSLVERR      (Logic0), 
           .PSEL         (PSEL), 
           .INTERRUPT    (INTERRUPT),
           .GP_OUT       (GP_OUT), 
           .GP_IN        (GP_IN), 
           .EXT_WR       (), 
           .EXT_RD       (), 
           .EXT_ADDR     (), 
           .EXT_DATA     (), 
           .EXT_WAIT     (Logic0), 
           .CON_ADDR     (), 
           .CON_DATA     (), 
           .CON_RD       (Logic0), 
           .CON_WR       (Logic0), 
           .CON_BUSY     (), 
           .FINISHED     (FINISHED), 
           .FAILED       (FAILED)
        );                       
                   
assign PRDATA = ( PSEL[1] ? PRDATA_1 : PRDATA_0) ;                   
                         
                         
/* #############################################################################
                         
SPIINT      Output interrupt 
SPISDO      Output serial data out (generated by SPI as master)
SPISS[7:0]  Output slave select (generated by SPI as master)
SPISCLKO    Output shift clock out (generated by SPI as master)
SPISDI      Input  shift data in (master or slave)
SPIRXAVAIL  Output request for data to be read - rx data available
SPITXRFM    Output indicates transmit done - ready for more
SPISSI      Input  slave select (when SPI in slave mode)
SPIOEN      Output output enable (when de-asserted output pad for SPISDO tri-stated). This is active when the SPI is writing output data and deactivated when there is not data to write. This signal is active high.
SPIMode     Output mode:  (when 1,  SPI is master, when 0, SPI is slave)

*/

// ********************************************************************************
// SPI Core - Master    

wire [7:0] M_SPISS;

CORESPI # (
  .APB_DWIDTH        (APB_DWIDTH),
  .CFG_FRAME_SIZE    (4),
  .FIFO_DEPTH        (4),
  .CFG_CLK           (2),
  .CFG_SPO           (1),
  .CFG_SPH           (1),
  .CFG_SPS           (0),
  .CFG_MODE          (0)
)USPIM ( //.TESTMODE   (1'b0),
                  .PCLK       (PCLK),   
                  .PRESETN    (PRESETN),
                  .PADDR      (PADDR[6:0]),  
                  .PSEL       (PSEL[0]),   
                  .PENABLE    (PENABLE),
                  .PWRITE     (PWRITE), 
                  .PWDATA     (PWDATA), 
                  .PRDATA    (PRDATA_0),

                  .SPISSI     (M_SPISSI), 
                  .SPISDI     (M_SPISDI), 
                  .SPICLKI    (M_SPICLKI),
                  .SPISS      (M_SPISS),  
                  .SPISCLKO   (M_SPISCLKO),  
                  .SPIOEN     (M_SPIOEN),    
                  .SPISDO     (M_SPISDO),    

                  .SPIINT     (GP_IN[0]), 
                  .SPIRXAVAIL (GP_IN[1]),
                  .SPITXRFM   (GP_IN[2]),  
                  .SPIMODE    (GP_IN[3]),
                  .PREADY     (),
                  .PSLVERR    ()

                  );

// ********************************************************************************
// SPI Core - Master    

wire [7:0] S_SPISS;


CORESPI # (
  .APB_DWIDTH        (APB_DWIDTH),
  .CFG_FRAME_SIZE    (4),
  .FIFO_DEPTH        (4),
  .CFG_CLK           (2),
  .CFG_SPO           (1),
  .CFG_SPH           (1),
  .CFG_SPS           (0),
  .CFG_MODE          (0)
)  USPIS ( //.TESTMODE   (1'b0),
                  .PCLK       (PCLK),   
                  .PRESETN    (PRESETN),
                  .PADDR      (PADDR[6:0]),  
                  .PSEL       (PSEL[1]),   
                  .PENABLE    (PENABLE),
                  .PWRITE     (PWRITE), 
                  .PWDATA     (PWDATA), 
                  .PRDATA    (PRDATA_1),

                  .SPISSI     (S_SPISSI), 
                  .SPISDI     (S_SPISDI), 
                  .SPICLKI    (S_SPICLKI),
                  .SPISS      (S_SPISS),  
                  .SPISCLKO   (S_SPISCLKO),  
                  .SPIOEN     (S_SPIOEN),    
                  .SPISDO     (S_SPISDO),    

                  .SPIINT     (GP_IN[8]), 
                  .SPIRXAVAIL (GP_IN[9]),
                  .SPITXRFM   (GP_IN[10]),  
                  .SPIMODE    (GP_IN[11]),
                  .PREADY     (),
                  .PSLVERR    ()

                  );



// *************************************************************************************
// SPI Connectivity

reg [31:0] shiftreg = 32'b000;

always @(posedge M_SPISCLKO)
begin
	shiftreg <= { shiftreg[30:0] , (M_SPISDO & M_SPIOEN)}; 
end

reg nscdata;
always @(negedge M_SPISCLKO)
begin
	nscdata <= shiftreg[8]; 
end
	

reg mux;
always @(*)
 begin
   case (GP_OUT[10:8])
     3'b000 :  mux = M_SPISDO & M_SPIOEN;
     3'b001 :  mux = M_SPISDO & M_SPIOEN;
     3'b010 :  mux = nscdata;			  // 9 clock delay
     3'b100 :  mux = S_SPISDO & S_SPIOEN;
     3'b101 :  mux = S_SPISDO & S_SPIOEN;
     3'b110 :  mux = S_SPISDO & S_SPIOEN;
	endcase
 end
 	
assign M_SPISDI  = mux;  
assign S_SPICLKI = M_SPISCLKO;
assign S_SPISSI  = M_SPISS[0];
assign S_SPISDI  = M_SPISDO & M_SPIOEN;


// For Waveform trace
wire SPICLK   =  M_SPISCLKO;
wire SPISEL   =  M_SPISS[0];
wire SPIDATAM =  M_SPISDO & M_SPIOEN;
wire SPIDATAS =  M_SPISDI;


// *************************************************************************************
// Simple Spy Capture Model

// AS: removed

//reg [7:0] capture = 8'b00;
//reg [7:0] capnext = 8'b00;
//integer bit = 0;

/*

always @(posedge SPICLK)
begin
  if (SPISEL==1)
  	 begin
  	   capture <= 8'b00;
      bit = 0;
    end 
  else
    begin
      capnext = { capture[6:0], M_SPISDO };
      capture <= capnext;
      bit = bit +1;
      if (bit==8)
       begin
       	$display("Captured %02d %02x",bit,capnext);
  	      capture <= 8'b00;
         bit = 0;
 		 end
 	 end	 	
end
    	  
*/

// *************************************************************************************
// PCLK Width Check

// AS: removed, not needed for USER TB

endmodule
