// ********************************************************************/
// Actel Corporation Proprietary and Confidential
// Copyright 2009 Actel Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
 //
//
// corespi.v
//
//
// Revision Information:
// Date     Description
//
//
// SVN Revision Information:
// SVN $Revision: 21608 $
// SVN $Date: 2013-12-02 16:03:36 -0800 (Mon, 02 Dec 2013) $
//
// Resolved SARs
// SAR      Date     Who   Description
// 72424       top level name
// 72425       PADDR 11 bits
// Notes:
//
//
// *********************************************************************/

module
CORESPI 
(	 //inputs
             PCLK,       //system clock
             PRESETN,    //system reset
             PADDR,      //address line
             PSEL,       //device select
             PENABLE,    //enable
             PWRITE,     //write
             PWDATA,     //write data
             SPISSI,     //slave select
             SPISDI,     //serial data in
             SPICLKI,    //serial clock in

             //outputs
             PRDATA,     //data read
             SPIINT,     //interrupt
             SPISS,      //slave select
             SPISCLKO,   //serial clock out
             SPIRXAVAIL, //data ready to be read (dma mode)
             SPITXRFM,   //room for more (dma mode)
             SPIOEN,     //output enable
             SPISDO,     //serial data out
             SPIMODE,     //1 -> master, 0 -> slave,
             PREADY,
             PSLVERR
             
             );

// AS: Added Parameters to replace 
// configuration bits / registers
parameter               FAMILY          =   15;
parameter               APB_DWIDTH      =   8;
parameter               CFG_FRAME_SIZE  =   4;
parameter               FIFO_DEPTH      =   4;
parameter               CFG_CLK         =   7;
parameter               CFG_SPO         =   0;
parameter               CFG_SPH         =   0;
parameter               CFG_SPS         =   0;
parameter               CFG_MODE        =   0;


//input TESTMODE;
input PCLK;
input PRESETN;
input [6:0] PADDR;
input PSEL;
input PENABLE;
input PWRITE;
input [APB_DWIDTH-1:0] PWDATA;
input SPISSI;
input SPISDI;
input SPICLKI;


output [APB_DWIDTH-1:0] PRDATA;
output SPIINT;
output [7:0] SPISS;
output SPISCLKO;
output SPIRXAVAIL;
output SPITXRFM;
output SPIOEN;
output SPIMODE;
output SPISDO;

// AP3
output PSLVERR;
output PREADY;

// tie off AP3 signals
assign PSLVERR = 1'b0;
assign PREADY = 1'b1;

spi # (
          .APB_DWIDTH     (APB_DWIDTH),
          .CFG_FRAME_SIZE (CFG_FRAME_SIZE),
          .FIFO_DEPTH     (FIFO_DEPTH),
          .CFG_CLK        (CFG_CLK),
          .CFG_SPO        (CFG_SPO),
          .CFG_SPH        (CFG_SPH),
          .CFG_SPS        (CFG_SPS),
          .CFG_MODE       (CFG_MODE)
) USPI( //inputs
//         .TESTMODE(TESTMODE),
         .PCLK(PCLK),      
         .PRESETN(PRESETN),
         .PADDR(PADDR),    
         .PSEL(PSEL),      
         .PENABLE(PENABLE),
         .PWRITE(PWRITE),  
         .PWDATA(PWDATA),  
         .SPISSI(SPISSI),  
         .SPISDI(SPISDI),  
         .SPICLKI(SPICLKI),
          
         //outputs
         .PRDDATA(PRDATA), 
         .SPIINT(SPIINT),  
         .SPISS(SPISS),    
         .SPISCLKO(SPISCLKO), 
         .SPIRXAVAIL(SPIRXAVAIL),
         .SPITXRFM(SPITXRFM), 
         .SPIOEN(SPIOEN), 
         .SPISDO(SPISDO), 
         .SPIMODE(SPIMODE)
         );

endmodule
